`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 02/12/2018 03:31:31 PM
// Design Name:
// Module Name: Font
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module FontROM(
	input wire [7:0] ascii,
	input wire [3:0] column,
	output wire [7:0] pixels
);

reg [7:0] out [0:16];
assign pixels = out[column];

always @(ascii or column) begin
	case(ascii)
		8'h00: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h01: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111110; // 2  ******
			out[3] <= 8'b10000001; // 3 *      *
			out[4] <= 8'b10100101; // 4 * *  * *
			out[5] <= 8'b10000001; // 5 *      *
			out[6] <= 8'b10000001; // 6 *      *
			out[7] <= 8'b10111101; // 7 * **** *
			out[8] <= 8'b10011001; // 8 *  **  *
			out[9] <= 8'b10000001; // 9 *      *
			out[10] <= 8'b10000001; // a *      *
			out[11] <= 8'b01111110; // b  ******
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h02: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111110; // 2  ******
			out[3] <= 8'b11111111; // 3 ********
			out[4] <= 8'b11011011; // 4 ** ** **
			out[5] <= 8'b11111111; // 5 ********
			out[6] <= 8'b11111111; // 6 ********
			out[7] <= 8'b11000011; // 7 **    **
			out[8] <= 8'b11100111; // 8 ***  ***
			out[9] <= 8'b11111111; // 9 ********
			out[10] <= 8'b11111111; // a ********
			out[11] <= 8'b01111110; // b  ******
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h03: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b01101100; // 4  ** **
			out[5] <= 8'b11111110; // 5 *******
			out[6] <= 8'b11111110; // 6 *******
			out[7] <= 8'b11111110; // 7 *******
			out[8] <= 8'b11111110; // 8 *******
			out[9] <= 8'b01111100; // 9  *****
			out[10] <= 8'b00111000; // a   ***
			out[11] <= 8'b00010000; // b    *
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h04: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00010000; // 4    *
			out[5] <= 8'b00111000; // 5   ***
			out[6] <= 8'b01111100; // 6  *****
			out[7] <= 8'b11111110; // 7 *******
			out[8] <= 8'b01111100; // 8  *****
			out[9] <= 8'b00111000; // 9   ***
			out[10] <= 8'b00010000; // a    *
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h05: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00011000; // 3    **
			out[4] <= 8'b00111100; // 4   ****
			out[5] <= 8'b00111100; // 5   ****
			out[6] <= 8'b11100111; // 6 ***  ***
			out[7] <= 8'b11100111; // 7 ***  ***
			out[8] <= 8'b11100111; // 8 ***  ***
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00111100; // b   ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h06: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00011000; // 3    **
			out[4] <= 8'b00111100; // 4   ****
			out[5] <= 8'b01111110; // 5  ******
			out[6] <= 8'b11111111; // 6 ********
			out[7] <= 8'b11111111; // 7 ********
			out[8] <= 8'b01111110; // 8  ******
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00111100; // b   ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h07: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00111100; // 7   ****
			out[8] <= 8'b00111100; // 8   ****
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		// 8'h08: begin
		// 	out[0] <= 8'b11111111; // 0 ********
		// 	out[1] <= 8'b11111111; // 1 ********
		// 	out[2] <= 8'b11111111; // 2 ********
		// 	out[3] <= 8'b11111111; // 3 ********
		// 	out[4] <= 8'b11111111; // 4 ********
		// 	out[5] <= 8'b11111111; // 5 ********
		// 	out[6] <= 8'b11100111; // 6 ***  ***
		// 	out[7] <= 8'b11000011; // 7 **    **
		// 	out[8] <= 8'b11000011; // 8 **    **
		// 	out[9] <= 8'b11100111; // 9 ***  ***
		// 	out[10] <= 8'b11111111; // a ********
		// 	out[11] <= 8'b11111111; // b ********
		// 	out[12] <= 8'b11111111; // c ********
		// 	out[13] <= 8'b11111111; // d ********
		// 	out[14] <= 8'b11111111; // e ********
		// 	out[15] <= 8'b11111111; // f ********
		// end
		"\n": begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h09: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00111100; // 5   ****
			out[6] <= 8'b01100110; // 6  **  **
			out[7] <= 8'b01000010; // 7  *    *
			out[8] <= 8'b01000010; // 8  *    *
			out[9] <= 8'b01100110; // 9  **  **
			out[10] <= 8'b00111100; // a   ****
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h0a: begin
			out[0] <= 8'b11111111; // 0 ********
			out[1] <= 8'b11111111; // 1 ********
			out[2] <= 8'b11111111; // 2 ********
			out[3] <= 8'b11111111; // 3 ********
			out[4] <= 8'b11111111; // 4 ********
			out[5] <= 8'b11000011; // 5 **    **
			out[6] <= 8'b10011001; // 6 *  **  *
			out[7] <= 8'b10111101; // 7 * **** *
			out[8] <= 8'b10111101; // 8 * **** *
			out[9] <= 8'b10011001; // 9 *  **  *
			out[10] <= 8'b11000011; // a **    **
			out[11] <= 8'b11111111; // b ********
			out[12] <= 8'b11111111; // c ********
			out[13] <= 8'b11111111; // d ********
			out[14] <= 8'b11111111; // e ********
			out[15] <= 8'b11111111; // f ********
		end
		8'h0b: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00011110; // 2    ****
			out[3] <= 8'b00001110; // 3     ***
			out[4] <= 8'b00011010; // 4    ** *
			out[5] <= 8'b00110010; // 5   **  *
			out[6] <= 8'b01111000; // 6  ****
			out[7] <= 8'b11001100; // 7 **  **
			out[8] <= 8'b11001100; // 8 **  **
			out[9] <= 8'b11001100; // 9 **  **
			out[10] <= 8'b11001100; // a **  **
			out[11] <= 8'b01111000; // b  ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h0c: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00111100; // 2   ****
			out[3] <= 8'b01100110; // 3  **  **
			out[4] <= 8'b01100110; // 4  **  **
			out[5] <= 8'b01100110; // 5  **  **
			out[6] <= 8'b01100110; // 6  **  **
			out[7] <= 8'b00111100; // 7   ****
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b01111110; // 9  ******
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00011000; // b    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h0d: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00111111; // 2   ******
			out[3] <= 8'b00110011; // 3   **  **
			out[4] <= 8'b00111111; // 4   ******
			out[5] <= 8'b00110000; // 5   **
			out[6] <= 8'b00110000; // 6   **
			out[7] <= 8'b00110000; // 7   **
			out[8] <= 8'b00110000; // 8   **
			out[9] <= 8'b01110000; // 9  ***
			out[10] <= 8'b11110000; // a ****
			out[11] <= 8'b11100000; // b ***
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h0e: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111111; // 2  *******
			out[3] <= 8'b01100011; // 3  **   **
			out[4] <= 8'b01111111; // 4  *******
			out[5] <= 8'b01100011; // 5  **   **
			out[6] <= 8'b01100011; // 6  **   **
			out[7] <= 8'b01100011; // 7  **   **
			out[8] <= 8'b01100011; // 8  **   **
			out[9] <= 8'b01100111; // 9  **  ***
			out[10] <= 8'b11100111; // a ***  ***
			out[11] <= 8'b11100110; // b ***  **
			out[12] <= 8'b11000000; // c **
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h0f: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00011000; // 3    **
			out[4] <= 8'b00011000; // 4    **
			out[5] <= 8'b11011011; // 5 ** ** **
			out[6] <= 8'b00111100; // 6   ****
			out[7] <= 8'b11100111; // 7 ***  ***
			out[8] <= 8'b00111100; // 8   ****
			out[9] <= 8'b11011011; // 9 ** ** **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00011000; // b    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h10: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b10000000; // 1 *
			out[2] <= 8'b11000000; // 2 **
			out[3] <= 8'b11100000; // 3 ***
			out[4] <= 8'b11110000; // 4 ****
			out[5] <= 8'b11111000; // 5 *****
			out[6] <= 8'b11111110; // 6 *******
			out[7] <= 8'b11111000; // 7 *****
			out[8] <= 8'b11110000; // 8 ****
			out[9] <= 8'b11100000; // 9 ***
			out[10] <= 8'b11000000; // a **
			out[11] <= 8'b10000000; // b *
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h11: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000010; // 1       *
			out[2] <= 8'b00000110; // 2      **
			out[3] <= 8'b00001110; // 3     ***
			out[4] <= 8'b00011110; // 4    ****
			out[5] <= 8'b00111110; // 5   *****
			out[6] <= 8'b11111110; // 6 *******
			out[7] <= 8'b00111110; // 7   *****
			out[8] <= 8'b00011110; // 8    ****
			out[9] <= 8'b00001110; // 9     ***
			out[10] <= 8'b00000110; // a      **
			out[11] <= 8'b00000010; // b       *
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h12: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00011000; // 2    **
			out[3] <= 8'b00111100; // 3   ****
			out[4] <= 8'b01111110; // 4  ******
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b01111110; // 8  ******
			out[9] <= 8'b00111100; // 9   ****
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h13: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01100110; // 2  **  **
			out[3] <= 8'b01100110; // 3  **  **
			out[4] <= 8'b01100110; // 4  **  **
			out[5] <= 8'b01100110; // 5  **  **
			out[6] <= 8'b01100110; // 6  **  **
			out[7] <= 8'b01100110; // 7  **  **
			out[8] <= 8'b01100110; // 8  **  **
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b01100110; // b  **  **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h14: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111111; // 2  *******
			out[3] <= 8'b11011011; // 3 ** ** **
			out[4] <= 8'b11011011; // 4 ** ** **
			out[5] <= 8'b11011011; // 5 ** ** **
			out[6] <= 8'b01111011; // 6  **** **
			out[7] <= 8'b00011011; // 7    ** **
			out[8] <= 8'b00011011; // 8    ** **
			out[9] <= 8'b00011011; // 9    ** **
			out[10] <= 8'b00011011; // a    ** **
			out[11] <= 8'b00011011; // b    ** **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h15: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b01111100; // 1  *****
			out[2] <= 8'b11000110; // 2 **   **
			out[3] <= 8'b01100000; // 3  **
			out[4] <= 8'b00111000; // 4   ***
			out[5] <= 8'b01101100; // 5  ** **
			out[6] <= 8'b11000110; // 6 **   **
			out[7] <= 8'b11000110; // 7 **   **
			out[8] <= 8'b01101100; // 8  ** **
			out[9] <= 8'b00111000; // 9   ***
			out[10] <= 8'b00001100; // a     **
			out[11] <= 8'b11000110; // b **   **
			out[12] <= 8'b01111100; // c  *****
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h16: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b11111110; // 8 *******
			out[9] <= 8'b11111110; // 9 *******
			out[10] <= 8'b11111110; // a *******
			out[11] <= 8'b11111110; // b *******
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h17: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00011000; // 2    **
			out[3] <= 8'b00111100; // 3   ****
			out[4] <= 8'b01111110; // 4  ******
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b01111110; // 8  ******
			out[9] <= 8'b00111100; // 9   ****
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b01111110; // b  ******
			out[12] <= 8'b00110000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h18: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00011000; // 2    **
			out[3] <= 8'b00111100; // 3   ****
			out[4] <= 8'b01111110; // 4  ******
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00011000; // b    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h19: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00011000; // 2    **
			out[3] <= 8'b00011000; // 3    **
			out[4] <= 8'b00011000; // 4    **
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b01111110; // 9  ******
			out[10] <= 8'b00111100; // a   ****
			out[11] <= 8'b00011000; // b    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h1a: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00001100; // 6     **
			out[7] <= 8'b11111110; // 7 *******
			out[8] <= 8'b00001100; // 8     **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h1b: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00110000; // 5   **
			out[6] <= 8'b01100000; // 6  **
			out[7] <= 8'b11111110; // 7 *******
			out[8] <= 8'b01100000; // 8  **
			out[9] <= 8'b00110000; // 9   **
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h1c: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b11000000; // 6 **
			out[7] <= 8'b11000000; // 7 **
			out[8] <= 8'b11000000; // 8 **
			out[9] <= 8'b11111110; // 9 *******
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h1d: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00100100; // 5   *  *
			out[6] <= 8'b01100110; // 6  **  **
			out[7] <= 8'b11111111; // 7 ********
			out[8] <= 8'b01100110; // 8  **  **
			out[9] <= 8'b00100100; // 9   *  *
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h1e: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00010000; // 4    *
			out[5] <= 8'b00111000; // 5   ***
			out[6] <= 8'b00111000; // 6   ***
			out[7] <= 8'b01111100; // 7  *****
			out[8] <= 8'b01111100; // 8  *****
			out[9] <= 8'b11111110; // 9 *******
			out[10] <= 8'b11111110; // a *******
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h1f: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b11111110; // 4 *******
			out[5] <= 8'b11111110; // 5 *******
			out[6] <= 8'b01111100; // 6  *****
			out[7] <= 8'b01111100; // 7  *****
			out[8] <= 8'b00111000; // 8   ***
			out[9] <= 8'b00111000; // 9   ***
			out[10] <= 8'b00010000; // a    *
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h20: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h21: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00011000; // 2    **
			out[3] <= 8'b00111100; // 3   ****
			out[4] <= 8'b00111100; // 4   ****
			out[5] <= 8'b00111100; // 5   ****
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00011000; // b    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h22: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b01100110; // 1  **  **
			out[2] <= 8'b01100110; // 2  **  **
			out[3] <= 8'b01100110; // 3  **  **
			out[4] <= 8'b00100100; // 4   *  *
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h23: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b01101100; // 3  ** **
			out[4] <= 8'b01101100; // 4  ** **
			out[5] <= 8'b11111110; // 5 *******
			out[6] <= 8'b01101100; // 6  ** **
			out[7] <= 8'b01101100; // 7  ** **
			out[8] <= 8'b01101100; // 8  ** **
			out[9] <= 8'b11111110; // 9 *******
			out[10] <= 8'b01101100; // a  ** **
			out[11] <= 8'b01101100; // b  ** **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h24: begin
			out[0] <= 8'b00011000; // 0     **
			out[1] <= 8'b00011000; // 1     **
			out[2] <= 8'b01111100; // 2   *****
			out[3] <= 8'b11000110; // 3  **   **
			out[4] <= 8'b11000010; // 4  **    *
			out[5] <= 8'b11000000; // 5  **
			out[6] <= 8'b01111100; // 6   *****
			out[7] <= 8'b00000110; // 7       **
			out[8] <= 8'b00000110; // 8       **
			out[9] <= 8'b10000110; // 9  *    **
			out[10] <= 8'b11000110; // a  **   **
			out[11] <= 8'b01111100; // b   *****
			out[12] <= 8'b00011000; // c     **
			out[13] <= 8'b00011000; // d     **
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h25: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b11000010; // 4 **    *
			out[5] <= 8'b11000110; // 5 **   **
			out[6] <= 8'b00001100; // 6     **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00110000; // 8   **
			out[9] <= 8'b01100000; // 9  **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b10000110; // b *    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h26: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00111000; // 2   ***
			out[3] <= 8'b01101100; // 3  ** **
			out[4] <= 8'b01101100; // 4  ** **
			out[5] <= 8'b00111000; // 5   ***
			out[6] <= 8'b01110110; // 6  *** **
			out[7] <= 8'b11011100; // 7 ** ***
			out[8] <= 8'b11001100; // 8 **  **
			out[9] <= 8'b11001100; // 9 **  **
			out[10] <= 8'b11001100; // a **  **
			out[11] <= 8'b01110110; // b  *** **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h27: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00110000; // 1   **
			out[2] <= 8'b00110000; // 2   **
			out[3] <= 8'b00110000; // 3   **
			out[4] <= 8'b01100000; // 4  **
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h28: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00001100; // 2     **
			out[3] <= 8'b00011000; // 3    **
			out[4] <= 8'b00110000; // 4   **
			out[5] <= 8'b00110000; // 5   **
			out[6] <= 8'b00110000; // 6   **
			out[7] <= 8'b00110000; // 7   **
			out[8] <= 8'b00110000; // 8   **
			out[9] <= 8'b00110000; // 9   **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00001100; // b     **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h29: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00110000; // 2   **
			out[3] <= 8'b00011000; // 3    **
			out[4] <= 8'b00001100; // 4     **
			out[5] <= 8'b00001100; // 5     **
			out[6] <= 8'b00001100; // 6     **
			out[7] <= 8'b00001100; // 7     **
			out[8] <= 8'b00001100; // 8     **
			out[9] <= 8'b00001100; // 9     **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00110000; // b   **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h2a: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b01100110; // 5  **  **
			out[6] <= 8'b00111100; // 6   ****
			out[7] <= 8'b11111111; // 7 ********
			out[8] <= 8'b00111100; // 8   ****
			out[9] <= 8'b01100110; // 9  **  **
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h2b: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b01111110; // 7  ******
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h2c: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00011000; // b    **
			out[12] <= 8'b00110000; // c   **
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h2d: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b01111110; // 7  ******
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h2e: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00011000; // b    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h2f: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000010; // 4       *
			out[5] <= 8'b00000110; // 5      **
			out[6] <= 8'b00001100; // 6     **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00110000; // 8   **
			out[9] <= 8'b01100000; // 9  **
			out[10] <= 8'b11000000; // a **
			out[11] <= 8'b10000000; // b *
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h30: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111100; // 2  *****
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b11000110; // 4 **   **
			out[5] <= 8'b11001110; // 5 **  ***
			out[6] <= 8'b11011110; // 6 ** ****
			out[7] <= 8'b11110110; // 7 **** **
			out[8] <= 8'b11100110; // 8 ***  **
			out[9] <= 8'b11000110; // 9 **   **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h31: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00011000; // 2
			out[3] <= 8'b00111000; // 3
			out[4] <= 8'b01111000; // 4    **
			out[5] <= 8'b00011000; // 5   ***
			out[6] <= 8'b00011000; // 6  ****
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b01111110; // b    **
			out[12] <= 8'b00000000; // c    **
			out[13] <= 8'b00000000; // d  ******
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h32: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111100; // 2  *****
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b00000110; // 4      **
			out[5] <= 8'b00001100; // 5     **
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00110000; // 7   **
			out[8] <= 8'b01100000; // 8  **
			out[9] <= 8'b11000000; // 9 **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b11111110; // b *******
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h33: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111100; // 2  *****
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b00000110; // 4      **
			out[5] <= 8'b00000110; // 5      **
			out[6] <= 8'b00111100; // 6   ****
			out[7] <= 8'b00000110; // 7      **
			out[8] <= 8'b00000110; // 8      **
			out[9] <= 8'b00000110; // 9      **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h34: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00001100; // 2     **
			out[3] <= 8'b00011100; // 3    ***
			out[4] <= 8'b00111100; // 4   ****
			out[5] <= 8'b01101100; // 5  ** **
			out[6] <= 8'b11001100; // 6 **  **
			out[7] <= 8'b11111110; // 7 *******
			out[8] <= 8'b00001100; // 8     **
			out[9] <= 8'b00001100; // 9     **
			out[10] <= 8'b00001100; // a     **
			out[11] <= 8'b00011110; // b    ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h35: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11111110; // 2 *******
			out[3] <= 8'b11000000; // 3 **
			out[4] <= 8'b11000000; // 4 **
			out[5] <= 8'b11000000; // 5 **
			out[6] <= 8'b11111100; // 6 ******
			out[7] <= 8'b00000110; // 7      **
			out[8] <= 8'b00000110; // 8      **
			out[9] <= 8'b00000110; // 9      **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h36: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00111000; // 2   ***
			out[3] <= 8'b01100000; // 3  **
			out[4] <= 8'b11000000; // 4 **
			out[5] <= 8'b11000000; // 5 **
			out[6] <= 8'b11111100; // 6 ******
			out[7] <= 8'b11000110; // 7 **   **
			out[8] <= 8'b11000110; // 8 **   **
			out[9] <= 8'b11000110; // 9 **   **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h37: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11111110; // 2 *******
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b00000110; // 4      **
			out[5] <= 8'b00000110; // 5      **
			out[6] <= 8'b00001100; // 6     **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00110000; // 8   **
			out[9] <= 8'b00110000; // 9   **
			out[10] <= 8'b00110000; // a   **
			out[11] <= 8'b00110000; // b   **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h38: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111100; // 2  *****
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b11000110; // 4 **   **
			out[5] <= 8'b11000110; // 5 **   **
			out[6] <= 8'b01111100; // 6  *****
			out[7] <= 8'b11000110; // 7 **   **
			out[8] <= 8'b11000110; // 8 **   **
			out[9] <= 8'b11000110; // 9 **   **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h39: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111100; // 2  *****
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b11000110; // 4 **   **
			out[5] <= 8'b11000110; // 5 **   **
			out[6] <= 8'b01111110; // 6  ******
			out[7] <= 8'b00000110; // 7      **
			out[8] <= 8'b00000110; // 8      **
			out[9] <= 8'b00000110; // 9      **
			out[10] <= 8'b00001100; // a     **
			out[11] <= 8'b01111000; // b  ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h3a: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00011000; // 4    **
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h3b: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00011000; // 4    **
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00110000; // b   **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h3c: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000110; // 3      **
			out[4] <= 8'b00001100; // 4     **
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00110000; // 6   **
			out[7] <= 8'b01100000; // 7  **
			out[8] <= 8'b00110000; // 8   **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00001100; // a     **
			out[11] <= 8'b00000110; // b      **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h3d: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b01111110; // 5  ******
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b01111110; // 8  ******
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h3e: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b01100000; // 3  **
			out[4] <= 8'b00110000; // 4   **
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00001100; // 6     **
			out[7] <= 8'b00000110; // 7      **
			out[8] <= 8'b00001100; // 8     **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00110000; // a   **
			out[11] <= 8'b01100000; // b  **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h3f: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111100; // 2  *****
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b11000110; // 4 **   **
			out[5] <= 8'b00001100; // 5     **
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00011000; // b    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h40: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111100; // 2  *****
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b11000110; // 4 **   **
			out[5] <= 8'b11000110; // 5 **   **
			out[6] <= 8'b11011110; // 6 ** ****
			out[7] <= 8'b11011110; // 7 ** ****
			out[8] <= 8'b11011110; // 8 ** ****
			out[9] <= 8'b11011100; // 9 ** ***
			out[10] <= 8'b11000000; // a **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h41: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00010000; // 2    *
			out[3] <= 8'b00111000; // 3   ***
			out[4] <= 8'b01101100; // 4  ** **
			out[5] <= 8'b11000110; // 5 **   **
			out[6] <= 8'b11000110; // 6 **   **
			out[7] <= 8'b11111110; // 7 *******
			out[8] <= 8'b11000110; // 8 **   **
			out[9] <= 8'b11000110; // 9 **   **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b11000110; // b **   **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h42: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11111100; // 2 ******
			out[3] <= 8'b01100110; // 3  **  **
			out[4] <= 8'b01100110; // 4  **  **
			out[5] <= 8'b01100110; // 5  **  **
			out[6] <= 8'b01111100; // 6  *****
			out[7] <= 8'b01100110; // 7  **  **
			out[8] <= 8'b01100110; // 8  **  **
			out[9] <= 8'b01100110; // 9  **  **
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b11111100; // b ******
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h43: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00111100; // 2   ****
			out[3] <= 8'b01100110; // 3  **  **
			out[4] <= 8'b11000010; // 4 **    *
			out[5] <= 8'b11000000; // 5 **
			out[6] <= 8'b11000000; // 6 **
			out[7] <= 8'b11000000; // 7 **
			out[8] <= 8'b11000000; // 8 **
			out[9] <= 8'b11000010; // 9 **    *
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b00111100; // b   ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h44: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11111000; // 2 *****
			out[3] <= 8'b01101100; // 3  ** **
			out[4] <= 8'b01100110; // 4  **  **
			out[5] <= 8'b01100110; // 5  **  **
			out[6] <= 8'b01100110; // 6  **  **
			out[7] <= 8'b01100110; // 7  **  **
			out[8] <= 8'b01100110; // 8  **  **
			out[9] <= 8'b01100110; // 9  **  **
			out[10] <= 8'b01101100; // a  ** **
			out[11] <= 8'b11111000; // b *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h45: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11111110; // 2 *******
			out[3] <= 8'b01100110; // 3  **  **
			out[4] <= 8'b01100010; // 4  **   *
			out[5] <= 8'b01101000; // 5  ** *
			out[6] <= 8'b01111000; // 6  ****
			out[7] <= 8'b01101000; // 7  ** *
			out[8] <= 8'b01100000; // 8  **
			out[9] <= 8'b01100010; // 9  **   *
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b11111110; // b *******
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h46: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11111110; // 2 *******
			out[3] <= 8'b01100110; // 3  **  **
			out[4] <= 8'b01100010; // 4  **   *
			out[5] <= 8'b01101000; // 5  ** *
			out[6] <= 8'b01111000; // 6  ****
			out[7] <= 8'b01101000; // 7  ** *
			out[8] <= 8'b01100000; // 8  **
			out[9] <= 8'b01100000; // 9  **
			out[10] <= 8'b01100000; // a  **
			out[11] <= 8'b11110000; // b ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h47: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00111100; // 2   ****
			out[3] <= 8'b01100110; // 3  **  **
			out[4] <= 8'b11000010; // 4 **    *
			out[5] <= 8'b11000000; // 5 **
			out[6] <= 8'b11000000; // 6 **
			out[7] <= 8'b11011110; // 7 ** ****
			out[8] <= 8'b11000110; // 8 **   **
			out[9] <= 8'b11000110; // 9 **   **
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b00111010; // b   *** *
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h48: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11000110; // 2 **   **
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b11000110; // 4 **   **
			out[5] <= 8'b11000110; // 5 **   **
			out[6] <= 8'b11111110; // 6 *******
			out[7] <= 8'b11000110; // 7 **   **
			out[8] <= 8'b11000110; // 8 **   **
			out[9] <= 8'b11000110; // 9 **   **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b11000110; // b **   **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h49: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00111100; // 2   ****
			out[3] <= 8'b00011000; // 3    **
			out[4] <= 8'b00011000; // 4    **
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00111100; // b   ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h4a: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00011110; // 2    ****
			out[3] <= 8'b00001100; // 3     **
			out[4] <= 8'b00001100; // 4     **
			out[5] <= 8'b00001100; // 5     **
			out[6] <= 8'b00001100; // 6     **
			out[7] <= 8'b00001100; // 7     **
			out[8] <= 8'b11001100; // 8 **  **
			out[9] <= 8'b11001100; // 9 **  **
			out[10] <= 8'b11001100; // a **  **
			out[11] <= 8'b01111000; // b  ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h4b: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11100110; // 2 ***  **
			out[3] <= 8'b01100110; // 3  **  **
			out[4] <= 8'b01100110; // 4  **  **
			out[5] <= 8'b01101100; // 5  ** **
			out[6] <= 8'b01111000; // 6  ****
			out[7] <= 8'b01111000; // 7  ****
			out[8] <= 8'b01101100; // 8  ** **
			out[9] <= 8'b01100110; // 9  **  **
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b11100110; // b ***  **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h4c: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11110000; // 2 ****
			out[3] <= 8'b01100000; // 3  **
			out[4] <= 8'b01100000; // 4  **
			out[5] <= 8'b01100000; // 5  **
			out[6] <= 8'b01100000; // 6  **
			out[7] <= 8'b01100000; // 7  **
			out[8] <= 8'b01100000; // 8  **
			out[9] <= 8'b01100010; // 9  **   *
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b11111110; // b *******
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h4d: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11000011; // 2 **    **
			out[3] <= 8'b11100111; // 3 ***  ***
			out[4] <= 8'b11111111; // 4 ********
			out[5] <= 8'b11111111; // 5 ********
			out[6] <= 8'b11011011; // 6 ** ** **
			out[7] <= 8'b11000011; // 7 **    **
			out[8] <= 8'b11000011; // 8 **    **
			out[9] <= 8'b11000011; // 9 **    **
			out[10] <= 8'b11000011; // a **    **
			out[11] <= 8'b11000011; // b **    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h4e: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11000110; // 2 **   **
			out[3] <= 8'b11100110; // 3 ***  **
			out[4] <= 8'b11110110; // 4 **** **
			out[5] <= 8'b11111110; // 5 *******
			out[6] <= 8'b11011110; // 6 ** ****
			out[7] <= 8'b11001110; // 7 **  ***
			out[8] <= 8'b11000110; // 8 **   **
			out[9] <= 8'b11000110; // 9 **   **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b11000110; // b **   **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h4f: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111100; // 2  *****
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b11000110; // 4 **   **
			out[5] <= 8'b11000110; // 5 **   **
			out[6] <= 8'b11000110; // 6 **   **
			out[7] <= 8'b11000110; // 7 **   **
			out[8] <= 8'b11000110; // 8 **   **
			out[9] <= 8'b11000110; // 9 **   **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h50: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11111100; // 2 ******
			out[3] <= 8'b01100110; // 3  **  **
			out[4] <= 8'b01100110; // 4  **  **
			out[5] <= 8'b01100110; // 5  **  **
			out[6] <= 8'b01111100; // 6  *****
			out[7] <= 8'b01100000; // 7  **
			out[8] <= 8'b01100000; // 8  **
			out[9] <= 8'b01100000; // 9  **
			out[10] <= 8'b01100000; // a  **
			out[11] <= 8'b11110000; // b ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h51: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111100; // 2  *****
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b11000110; // 4 **   **
			out[5] <= 8'b11000110; // 5 **   **
			out[6] <= 8'b11000110; // 6 **   **
			out[7] <= 8'b11000110; // 7 **   **
			out[8] <= 8'b11000110; // 8 **   **
			out[9] <= 8'b11010110; // 9 ** * **
			out[10] <= 8'b11011110; // a ** ****
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00001100; // c     **
			out[13] <= 8'b00001110; // d     ***
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h52: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11111100; // 2 ******
			out[3] <= 8'b01100110; // 3  **  **
			out[4] <= 8'b01100110; // 4  **  **
			out[5] <= 8'b01100110; // 5  **  **
			out[6] <= 8'b01111100; // 6  *****
			out[7] <= 8'b01101100; // 7  ** **
			out[8] <= 8'b01100110; // 8  **  **
			out[9] <= 8'b01100110; // 9  **  **
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b11100110; // b ***  **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h53: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01111100; // 2  *****
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b11000110; // 4 **   **
			out[5] <= 8'b01100000; // 5  **
			out[6] <= 8'b00111000; // 6   ***
			out[7] <= 8'b00001100; // 7     **
			out[8] <= 8'b00000110; // 8      **
			out[9] <= 8'b11000110; // 9 **   **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h54: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11111111; // 2 ********
			out[3] <= 8'b11011011; // 3 ** ** **
			out[4] <= 8'b10011001; // 4 *  **  *
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00111100; // b   ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h55: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11000110; // 2 **   **
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b11000110; // 4 **   **
			out[5] <= 8'b11000110; // 5 **   **
			out[6] <= 8'b11000110; // 6 **   **
			out[7] <= 8'b11000110; // 7 **   **
			out[8] <= 8'b11000110; // 8 **   **
			out[9] <= 8'b11000110; // 9 **   **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h56: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11000011; // 2 **    **
			out[3] <= 8'b11000011; // 3 **    **
			out[4] <= 8'b11000011; // 4 **    **
			out[5] <= 8'b11000011; // 5 **    **
			out[6] <= 8'b11000011; // 6 **    **
			out[7] <= 8'b11000011; // 7 **    **
			out[8] <= 8'b11000011; // 8 **    **
			out[9] <= 8'b01100110; // 9  **  **
			out[10] <= 8'b00111100; // a   ****
			out[11] <= 8'b00011000; // b    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h57: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11000011; // 2 **    **
			out[3] <= 8'b11000011; // 3 **    **
			out[4] <= 8'b11000011; // 4 **    **
			out[5] <= 8'b11000011; // 5 **    **
			out[6] <= 8'b11000011; // 6 **    **
			out[7] <= 8'b11011011; // 7 ** ** **
			out[8] <= 8'b11011011; // 8 ** ** **
			out[9] <= 8'b11111111; // 9 ********
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b01100110; // b  **  **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h58: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11000011; // 2 **    **
			out[3] <= 8'b11000011; // 3 **    **
			out[4] <= 8'b01100110; // 4  **  **
			out[5] <= 8'b00111100; // 5   ****
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00111100; // 8   ****
			out[9] <= 8'b01100110; // 9  **  **
			out[10] <= 8'b11000011; // a **    **
			out[11] <= 8'b11000011; // b **    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h59: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11000011; // 2 **    **
			out[3] <= 8'b11000011; // 3 **    **
			out[4] <= 8'b11000011; // 4 **    **
			out[5] <= 8'b01100110; // 5  **  **
			out[6] <= 8'b00111100; // 6   ****
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00111100; // b   ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h5a: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11111111; // 2 ********
			out[3] <= 8'b11000011; // 3 **    **
			out[4] <= 8'b10000110; // 4 *    **
			out[5] <= 8'b00001100; // 5     **
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00110000; // 7   **
			out[8] <= 8'b01100000; // 8  **
			out[9] <= 8'b11000001; // 9 **     *
			out[10] <= 8'b11000011; // a **    **
			out[11] <= 8'b11111111; // b ********
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h5b: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00111100; // 2   ****
			out[3] <= 8'b00110000; // 3   **
			out[4] <= 8'b00110000; // 4   **
			out[5] <= 8'b00110000; // 5   **
			out[6] <= 8'b00110000; // 6   **
			out[7] <= 8'b00110000; // 7   **
			out[8] <= 8'b00110000; // 8   **
			out[9] <= 8'b00110000; // 9   **
			out[10] <= 8'b00110000; // a   **
			out[11] <= 8'b00111100; // b   ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h5c: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b10000000; // 3 *
			out[4] <= 8'b11000000; // 4 **
			out[5] <= 8'b11100000; // 5 ***
			out[6] <= 8'b01110000; // 6  ***
			out[7] <= 8'b00111000; // 7   ***
			out[8] <= 8'b00011100; // 8    ***
			out[9] <= 8'b00001110; // 9     ***
			out[10] <= 8'b00000110; // a      **
			out[11] <= 8'b00000010; // b       *
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h5d: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00111100; // 2   ****
			out[3] <= 8'b00001100; // 3     **
			out[4] <= 8'b00001100; // 4     **
			out[5] <= 8'b00001100; // 5     **
			out[6] <= 8'b00001100; // 6     **
			out[7] <= 8'b00001100; // 7     **
			out[8] <= 8'b00001100; // 8     **
			out[9] <= 8'b00001100; // 9     **
			out[10] <= 8'b00001100; // a     **
			out[11] <= 8'b00111100; // b   ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h5e: begin
			out[0] <= 8'b00010000; // 0    *
			out[1] <= 8'b00111000; // 1   ***
			out[2] <= 8'b01101100; // 2  ** **
			out[3] <= 8'b11000110; // 3 **   **
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h5f: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b11111111; // d ********
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h60: begin
			out[0] <= 8'b00110000; // 0   **
			out[1] <= 8'b00110000; // 1   **
			out[2] <= 8'b00011000; // 2    **
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h61: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b01111000; // 5  ****
			out[6] <= 8'b00001100; // 6     **
			out[7] <= 8'b01111100; // 7  *****
			out[8] <= 8'b11001100; // 8 **  **
			out[9] <= 8'b11001100; // 9 **  **
			out[10] <= 8'b11001100; // a **  **
			out[11] <= 8'b01110110; // b  *** **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h62: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11100000; // 2  ***
			out[3] <= 8'b01100000; // 3   **
			out[4] <= 8'b01100000; // 4   **
			out[5] <= 8'b01111000; // 5   ****
			out[6] <= 8'b01101100; // 6   ** **
			out[7] <= 8'b01100110; // 7   **  **
			out[8] <= 8'b01100110; // 8   **  **
			out[9] <= 8'b01100110; // 9   **  **
			out[10] <= 8'b01100110; // a   **  **
			out[11] <= 8'b01111100; // b   *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h63: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b01111100; // 5  *****
			out[6] <= 8'b11000110; // 6 **   **
			out[7] <= 8'b11000000; // 7 **
			out[8] <= 8'b11000000; // 8 **
			out[9] <= 8'b11000000; // 9 **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h64: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00011100; // 2    ***
			out[3] <= 8'b00001100; // 3     **
			out[4] <= 8'b00001100; // 4     **
			out[5] <= 8'b00111100; // 5   ****
			out[6] <= 8'b01101100; // 6  ** **
			out[7] <= 8'b11001100; // 7 **  **
			out[8] <= 8'b11001100; // 8 **  **
			out[9] <= 8'b11001100; // 9 **  **
			out[10] <= 8'b11001100; // a **  **
			out[11] <= 8'b01110110; // b  *** **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h65: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b01111100; // 5  *****
			out[6] <= 8'b11000110; // 6 **   **
			out[7] <= 8'b11111110; // 7 *******
			out[8] <= 8'b11000000; // 8 **
			out[9] <= 8'b11000000; // 9 **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h66: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00111000; // 2   ***
			out[3] <= 8'b01101100; // 3  ** **
			out[4] <= 8'b01100100; // 4  **  *
			out[5] <= 8'b01100000; // 5  **
			out[6] <= 8'b11110000; // 6 ****
			out[7] <= 8'b01100000; // 7  **
			out[8] <= 8'b01100000; // 8  **
			out[9] <= 8'b01100000; // 9  **
			out[10] <= 8'b01100000; // a  **
			out[11] <= 8'b11110000; // b ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h67: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b01110110; // 5  *** **
			out[6] <= 8'b11001100; // 6 **  **
			out[7] <= 8'b11001100; // 7 **  **
			out[8] <= 8'b11001100; // 8 **  **
			out[9] <= 8'b11001100; // 9 **  **
			out[10] <= 8'b11001100; // a **  **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00001100; // c     **
			out[13] <= 8'b11001100; // d **  **
			out[14] <= 8'b01111000; // e  ****
			out[15] <= 8'b00000000; // f
		end
		8'h68: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11100000; // 2 ***
			out[3] <= 8'b01100000; // 3  **
			out[4] <= 8'b01100000; // 4  **
			out[5] <= 8'b01101100; // 5  ** **
			out[6] <= 8'b01110110; // 6  *** **
			out[7] <= 8'b01100110; // 7  **  **
			out[8] <= 8'b01100110; // 8  **  **
			out[9] <= 8'b01100110; // 9  **  **
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b11100110; // b ***  **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h69: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00011000; // 2    **
			out[3] <= 8'b00011000; // 3    **
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00111000; // 5   ***
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00111100; // b   ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h6a: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000110; // 2      **
			out[3] <= 8'b00000110; // 3      **
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00001110; // 5     ***
			out[6] <= 8'b00000110; // 6      **
			out[7] <= 8'b00000110; // 7      **
			out[8] <= 8'b00000110; // 8      **
			out[9] <= 8'b00000110; // 9      **
			out[10] <= 8'b00000110; // a      **
			out[11] <= 8'b00000110; // b      **
			out[12] <= 8'b01100110; // c  **  **
			out[13] <= 8'b01100110; // d  **  **
			out[14] <= 8'b00111100; // e   ****
			out[15] <= 8'b00000000; // f
		end
		8'h6b: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b11100000; // 2 ***
			out[3] <= 8'b01100000; // 3  **
			out[4] <= 8'b01100000; // 4  **
			out[5] <= 8'b01100110; // 5  **  **
			out[6] <= 8'b01101100; // 6  ** **
			out[7] <= 8'b01111000; // 7  ****
			out[8] <= 8'b01111000; // 8  ****
			out[9] <= 8'b01101100; // 9  ** **
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b11100110; // b ***  **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h6c: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00111000; // 2   ***
			out[3] <= 8'b00011000; // 3    **
			out[4] <= 8'b00011000; // 4    **
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00011000; // 6    **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00111100; // b   ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h6d: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b11100110; // 5 ***  **
			out[6] <= 8'b11111111; // 6 ********
			out[7] <= 8'b11011011; // 7 ** ** **
			out[8] <= 8'b11011011; // 8 ** ** **
			out[9] <= 8'b11011011; // 9 ** ** **
			out[10] <= 8'b11011011; // a ** ** **
			out[11] <= 8'b11011011; // b ** ** **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h6e: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b11011100; // 5 ** ***
			out[6] <= 8'b01100110; // 6  **  **
			out[7] <= 8'b01100110; // 7  **  **
			out[8] <= 8'b01100110; // 8  **  **
			out[9] <= 8'b01100110; // 9  **  **
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b01100110; // b  **  **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h6f: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b01111100; // 5  *****
			out[6] <= 8'b11000110; // 6 **   **
			out[7] <= 8'b11000110; // 7 **   **
			out[8] <= 8'b11000110; // 8 **   **
			out[9] <= 8'b11000110; // 9 **   **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h70: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b11011100; // 5 ** ***
			out[6] <= 8'b01100110; // 6  **  **
			out[7] <= 8'b01100110; // 7  **  **
			out[8] <= 8'b01100110; // 8  **  **
			out[9] <= 8'b01100110; // 9  **  **
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b01100000; // c  **
			out[13] <= 8'b01100000; // d  **
			out[14] <= 8'b11110000; // e ****
			out[15] <= 8'b00000000; // f
		end
		8'h71: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b01110110; // 5  *** **
			out[6] <= 8'b11001100; // 6 **  **
			out[7] <= 8'b11001100; // 7 **  **
			out[8] <= 8'b11001100; // 8 **  **
			out[9] <= 8'b11001100; // 9 **  **
			out[10] <= 8'b11001100; // a **  **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00001100; // c     **
			out[13] <= 8'b00001100; // d     **
			out[14] <= 8'b00011110; // e    ****
			out[15] <= 8'b00000000; // f
		end
		8'h72: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b11011100; // 5 ** ***
			out[6] <= 8'b01110110; // 6  *** **
			out[7] <= 8'b01100110; // 7  **  **
			out[8] <= 8'b01100000; // 8  **
			out[9] <= 8'b01100000; // 9  **
			out[10] <= 8'b01100000; // a  **
			out[11] <= 8'b11110000; // b ****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h73: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b01111100; // 5  *****
			out[6] <= 8'b11000110; // 6 **   **
			out[7] <= 8'b01100000; // 7  **
			out[8] <= 8'b00111000; // 8   ***
			out[9] <= 8'b00001100; // 9     **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b01111100; // b  *****
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h74: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00010000; // 2    *
			out[3] <= 8'b00110000; // 3   **
			out[4] <= 8'b00110000; // 4   **
			out[5] <= 8'b11111100; // 5 ******
			out[6] <= 8'b00110000; // 6   **
			out[7] <= 8'b00110000; // 7   **
			out[8] <= 8'b00110000; // 8   **
			out[9] <= 8'b00110000; // 9   **
			out[10] <= 8'b00110110; // a   ** **
			out[11] <= 8'b00011100; // b    ***
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h75: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b11001100; // 5 **  **
			out[6] <= 8'b11001100; // 6 **  **
			out[7] <= 8'b11001100; // 7 **  **
			out[8] <= 8'b11001100; // 8 **  **
			out[9] <= 8'b11001100; // 9 **  **
			out[10] <= 8'b11001100; // a **  **
			out[11] <= 8'b01110110; // b  *** **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h76: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b11000011; // 5 **    **
			out[6] <= 8'b11000011; // 6 **    **
			out[7] <= 8'b11000011; // 7 **    **
			out[8] <= 8'b11000011; // 8 **    **
			out[9] <= 8'b01100110; // 9  **  **
			out[10] <= 8'b00111100; // a   ****
			out[11] <= 8'b00011000; // b    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h77: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b11000011; // 5 **    **
			out[6] <= 8'b11000011; // 6 **    **
			out[7] <= 8'b11000011; // 7 **    **
			out[8] <= 8'b11011011; // 8 ** ** **
			out[9] <= 8'b11011011; // 9 ** ** **
			out[10] <= 8'b11111111; // a ********
			out[11] <= 8'b01100110; // b  **  **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h78: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b11000011; // 5 **    **
			out[6] <= 8'b01100110; // 6  **  **
			out[7] <= 8'b00111100; // 7   ****
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00111100; // 9   ****
			out[10] <= 8'b01100110; // a  **  **
			out[11] <= 8'b11000011; // b **    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h79: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b11000110; // 5 **   **
			out[6] <= 8'b11000110; // 6 **   **
			out[7] <= 8'b11000110; // 7 **   **
			out[8] <= 8'b11000110; // 8 **   **
			out[9] <= 8'b11000110; // 9 **   **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b01111110; // b  ******
			out[12] <= 8'b00000110; // c      **
			out[13] <= 8'b00001100; // d     **
			out[14] <= 8'b11111000; // e *****
			out[15] <= 8'b00000000; // f
		end
		8'h7a: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b11111110; // 5 *******
			out[6] <= 8'b11001100; // 6 **  **
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00110000; // 8   **
			out[9] <= 8'b01100000; // 9  **
			out[10] <= 8'b11000110; // a **   **
			out[11] <= 8'b11111110; // b *******
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h7b: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00001110; // 2     ***
			out[3] <= 8'b00011000; // 3    **
			out[4] <= 8'b00011000; // 4    **
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b01110000; // 6  ***
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00001110; // b     ***
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h7c: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00011000; // 2    **
			out[3] <= 8'b00011000; // 3    **
			out[4] <= 8'b00011000; // 4    **
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b00011000; // b    **
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h7d: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01110000; // 2  ***
			out[3] <= 8'b00011000; // 3    **
			out[4] <= 8'b00011000; // 4    **
			out[5] <= 8'b00011000; // 5    **
			out[6] <= 8'b00001110; // 6     ***
			out[7] <= 8'b00011000; // 7    **
			out[8] <= 8'b00011000; // 8    **
			out[9] <= 8'b00011000; // 9    **
			out[10] <= 8'b00011000; // a    **
			out[11] <= 8'b01110000; // b  ***
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h7e: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b01110110; // 2  *** **
			out[3] <= 8'b11011100; // 3 ** ***
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000; // f
		end
		8'h7f: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00010000; // 4    *
			out[5] <= 8'b00111000; // 5   ***
			out[6] <= 8'b01101100; // 6  ** **
			out[7] <= 8'b11000110; // 7 **   **
			out[8] <= 8'b11000110; // 8 **   **
			out[9] <= 8'b11000110; // 9 **   **
			out[10] <= 8'b11111110; // a *******
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000;  // f
		end
		8'h80: begin
			out[0] <= 8'b11111111; // 0 ********
			out[1] <= 8'b11111111; // 1 ********
			out[2] <= 8'b11111111; // 2 ********
			out[3] <= 8'b11111111; // 3 ********
			out[4] <= 8'b11111111; // 4 ********
			out[5] <= 8'b11111111; // 5 ********
			out[6] <= 8'b11100111; // 6 ***  ***
			out[7] <= 8'b11000011; // 7 **    **
			out[8] <= 8'b11000011; // 8 **    **
			out[9] <= 8'b11100111; // 9 ***  ***
			out[10] <= 8'b11111111; // a ********
			out[11] <= 8'b11111111; // b ********
			out[12] <= 8'b11111111; // c ********
			out[13] <= 8'b11111111; // d ********
			out[14] <= 8'b11111111; // e ********
			out[15] <= 8'b11111111; // f ********
		end
		8'h81: begin
			out[0] <= 8'b11111111; // 0 ********
			out[1] <= 8'b11111111; // 1 ********
			out[2] <= 8'b11111111; // 2 ********
			out[3] <= 8'b11111111; // 3 ********
			out[4] <= 8'b11111111; // 4 ********
			out[5] <= 8'b11111111; // 5 ********
			out[6] <= 8'b11111111; // 6 ********
			out[7] <= 8'b11111111; // 7 ********
			out[8] <= 8'b11111111; // 8 ********
			out[9] <= 8'b11111111; // 9 ********
			out[10] <= 8'b11111111; // a ********
			out[11] <= 8'b11111111; // b ********
			out[12] <= 8'b11111111; // c ********
			out[13] <= 8'b11111111; // d ********
			out[14] <= 8'b11111111; // e ********
			out[15] <= 8'b11111111; // f ********
		end
		default: begin
			out[0] <= 8'b00000000; // 0
			out[1] <= 8'b00000000; // 1
			out[2] <= 8'b00000000; // 2
			out[3] <= 8'b00000000; // 3
			out[4] <= 8'b00000000; // 4
			out[5] <= 8'b00000000; // 5
			out[6] <= 8'b00000000; // 6
			out[7] <= 8'b00000000; // 7
			out[8] <= 8'b00000000; // 8
			out[9] <= 8'b00000000; // 9
			out[10] <= 8'b00000000; // a
			out[11] <= 8'b00000000; // b
			out[12] <= 8'b00000000; // c
			out[13] <= 8'b00000000; // d
			out[14] <= 8'b00000000; // e
			out[15] <= 8'b00000000;  // f
		end
	endcase
end
endmodule